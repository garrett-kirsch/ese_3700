*** SPICE deck for cell not{sch} from library ese3700
*** Created on Thu Feb 20, 2025 17:47:38
*** Last revised on Thu Feb 20, 2025 17:49:17
*** Written on Thu Feb 20, 2025 17:52:28 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: not{sch}
Mnmos@0 net@0 net@2 gnd gnd N L=0.022U W=0.044U
Mpmos@0 vdd net@2 net@0 vdd P L=0.022U W=0.044U
VV_Generi@0 vdd gnd DC 0.5 AC 0
VV_Generi@1 net@2 gnd DC 0 AC 0
.END
