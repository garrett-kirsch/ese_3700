*** SPICE deck for cell hw3_3b{sch} from library ese3700
*** Created on Wed Feb 12, 2025 16:24:30
*** Last revised on Wed Feb 12, 2025 16:32:57
*** Written on Wed Feb 12, 2025 16:33:14 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: hw3_3b{sch}
Mnmos@0 net@20 net@6 gnd gnd N L=0.022U W=0.022U
Mnmos@1 vdd net@20 gnd gnd N L=0.022U W=0.022U
Mnmos@2 vdd net@20 gnd gnd N L=0.022U W=0.022U
Mnmos@3 vdd net@20 gnd gnd N L=0.022U W=0.022U
Mnmos@4 vdd net@20 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@6 net@20 vdd P L=0.022U W=0.022U
VVPulse@0 net@6 gnd pulse (0.8V 0V 0ns 2ps 2ps 3ns 6ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
.END
