*** SPICE deck for cell test_single_sram{sch} from library ese_3700_project_2
*** Created on Fri May 02, 2025 13:59:51
*** Last revised on Fri May 02, 2025 23:12:00
*** Written on Fri May 02, 2025 23:12:06 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

*** SUBCIRCUIT ese_3700_project_2__not FROM CELL not{sch}
.SUBCKT ese_3700_project_2__not IN OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd IN OUT vdd P L=0.022U W=0.022U
.ENDS ese_3700_project_2__not

*** SUBCIRCUIT ese_3700_project_2__SRAM_CELL FROM CELL SRAM_CELL{sch}
.SUBCKT ese_3700_project_2__SRAM_CELL /BL BL WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 WL BL gnd N L=0.022U W=0.022U
Mnmos@1 /BL WL net@3 gnd N L=0.022U W=0.022U
Xnot@0 net@0 net@3 ese_3700_project_2__not
Xnot@1 net@3 net@0 ese_3700_project_2__not
.ENDS ese_3700_project_2__SRAM_CELL

*** SUBCIRCUIT ese_3700_project_2__nand2 FROM CELL nand2{sch}
.SUBCKT ese_3700_project_2__nand2 A B OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT A net@1 gnd N L=0.022U W=0.022U
Mnmos@1 net@1 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A OUT vdd P L=0.022U W=0.022U
Mpmos@1 vdd B OUT vdd P L=0.022U W=0.022U
.ENDS ese_3700_project_2__nand2

*** SUBCIRCUIT ese_3700_project_2__read_precharger FROM CELL read_precharger{sch}
.SUBCKT ese_3700_project_2__read_precharger _BL _Pre BL
** GLOBAL vdd
Mpmos@0 vdd _Pre BL vdd P L=0.022U W=0.176U
Mpmos@1 vdd _Pre _BL vdd P L=0.022U W=0.176U
Mpmos@2 BL _Pre _BL vdd P L=0.022U W=0.176U
.ENDS ese_3700_project_2__read_precharger

*** SUBCIRCUIT ese_3700_project_2__latch FROM CELL latch{sch}
.SUBCKT ese_3700_project_2__latch CLK IN OUT
** GLOBAL gnd
** GLOBAL vdd
Xnand2@3 IN CLK net@29 ese_3700_project_2__nand2
Xnand2@4 net@26 OUT net@27 ese_3700_project_2__nand2
Xnand2@5 net@29 net@27 OUT ese_3700_project_2__nand2
Xnot@1 CLK net@26 ese_3700_project_2__not
.ENDS ese_3700_project_2__latch

*** SUBCIRCUIT ese_3700_project_2__register FROM CELL register{sch}
.SUBCKT ese_3700_project_2__register _CLK CLK IN OUT
** GLOBAL gnd
** GLOBAL vdd
Xlatch@2 _CLK IN net@19 ese_3700_project_2__latch
Xlatch@3 CLK net@19 OUT ese_3700_project_2__latch
.ENDS ese_3700_project_2__register

*** SUBCIRCUIT ese_3700_project_2__tristate_buffer FROM CELL tristate_buffer{sch}
.SUBCKT ese_3700_project_2__tristate_buffer Enable In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@22 In gnd gnd N L=0.022U W=0.022U
Mnmos@1 out Enable net@28 gnd N L=0.022U W=0.022U
Mnmos@2 net@28 net@22 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@34 Enable gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd In net@22 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@22 net@26 vdd P L=0.022U W=0.022U
Mpmos@2 net@26 net@34 out vdd P L=0.022U W=0.022U
Mpmos@3 vdd Enable net@34 vdd P L=0.022U W=0.022U
.ENDS ese_3700_project_2__tristate_buffer

*** SUBCIRCUIT ese_3700_project_2__tristate_enable_inverter FROM CELL tristate_enable_inverter{sch}
.SUBCKT ese_3700_project_2__tristate_enable_inverter Enable In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@22 In gnd gnd N L=0.022U W=0.022U
Mnmos@1 out net@34 net@28 gnd N L=0.022U W=0.022U
Mnmos@2 net@28 net@22 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@34 Enable gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd In net@22 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@22 net@26 vdd P L=0.022U W=0.022U
Mpmos@2 net@26 Enable out vdd P L=0.022U W=0.022U
Mpmos@3 vdd Enable net@34 vdd P L=0.022U W=0.022U
.ENDS ese_3700_project_2__tristate_enable_inverter

*** SUBCIRCUIT ese_3700_project_2__tristate_driver FROM CELL tristate_driver{sch}
.SUBCKT ese_3700_project_2__tristate_driver _rd/wr BL cs d_in d_out
** GLOBAL gnd
** GLOBAL vdd
Xtristate@1 _rd/wr net@0 BL ese_3700_project_2__tristate_buffer
Xtristate@3 cs net@3 d_out ese_3700_project_2__tristate_buffer
Xtristate@4 cs d_in net@0 ese_3700_project_2__tristate_buffer
Xtristate@6 _rd/wr BL net@3 ese_3700_project_2__tristate_enable_inverter
.ENDS ese_3700_project_2__tristate_driver

*** SUBCIRCUIT ese_3700_project_2__tristate_inverter FROM CELL tristate_inverter{sch}
.SUBCKT ese_3700_project_2__tristate_inverter Enable In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 out Enable net@28 gnd N L=0.022U W=0.022U
Mnmos@2 net@28 In gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@34 Enable gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd In net@26 vdd P L=0.022U W=0.022U
Mpmos@2 net@26 net@34 out vdd P L=0.022U W=0.022U
Mpmos@3 vdd Enable net@34 vdd P L=0.022U W=0.022U
.ENDS ese_3700_project_2__tristate_inverter

*** SUBCIRCUIT hw6__buffer FROM CELL hw6:buffer{sch}
.SUBCKT hw6__buffer IN OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@26 IN gnd gnd N L=0.022U W=0.022U
Mnmos@2 OUT net@26 gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd IN net@26 vdd P L=0.022U W=0.022U
Mpmos@2 vdd net@26 OUT vdd P L=0.022U W=0.022U
.ENDS hw6__buffer

*** SUBCIRCUIT hw6__nor2 FROM CELL hw6:nor2{sch}
.SUBCKT hw6__nor2 A B OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT A gnd gnd N L=0.022U W=0.022U
Mnmos@1 OUT B gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@2 B OUT vdd P L=0.022U W=0.022U
Mpmos@1 vdd A net@2 vdd P L=0.022U W=0.022U
.ENDS hw6__nor2

*** SUBCIRCUIT ese_3700_project_2__two_phase_clock_generator FROM CELL two_phase_clock_generator{sch}
.SUBCKT ese_3700_project_2__two_phase_clock_generator _CLK CLK IN
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 IN b hw6__buffer
Xnor2@0 a _CLK CLK hw6__nor2
Xnor2@1 CLK b _CLK hw6__nor2
Xnot@0 IN a ese_3700_project_2__not
.ENDS ese_3700_project_2__two_phase_clock_generator

*** SUBCIRCUIT ese_3700_project_2__single_cell_sram FROM CELL single_cell_sram{sch}
.SUBCKT ese_3700_project_2__single_cell_sram _rd/wr CLK_in d_in d_out
** GLOBAL gnd
** GLOBAL vdd
XSRAM_CEL@0 net@35 net@12 net@43 ese_3700_project_2__SRAM_CELL
Xnand2@0 net@41 net@54 net@57 ese_3700_project_2__nand2
Xnot@0 net@4 net@54 ese_3700_project_2__not
Xread_pre@0 net@35 net@57 net@12 ese_3700_project_2__read_precharger
Xregister@0 net@43 net@41 _rd/wr net@4 ese_3700_project_2__register
Xregister@1 net@43 net@41 d_in net@19 ese_3700_project_2__register
Xregister@2 net@43 net@41 net@71 d_out ese_3700_project_2__register
Xtristate@0 net@4 net@12 vdd net@19 net@71 ese_3700_project_2__tristate_driver
Xtristate@5 net@4 net@12 net@35 ese_3700_project_2__tristate_inverter
Xtwo_phas@0 net@43 net@41 CLK_in ese_3700_project_2__two_phase_clock_generator
.ENDS ese_3700_project_2__single_cell_sram

.global gnd vdd

*** TOP LEVEL CELL: test_single_sram{sch}
VVPWL@0 wr gnd pulse (0V 0.8V 0ns 1ps 1ps 2ns 6ns) DC 0V AC 0V 0
VVPulse@0 CLK gnd pulse (0.8V 0V 0ns 1ps 1ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@1 din gnd pulse (0V 0.8V 0ns 1ps 1ps 12ns 24ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xsingle_c@0 wr CLK din dout ese_3700_project_2__single_cell_sram
.END
