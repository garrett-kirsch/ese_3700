*** SPICE deck for cell hw2_tranisient{sch} from library ese3700
*** Created on Sat Feb 08, 2025 11:42:36
*** Last revised on Sat Feb 08, 2025 12:56:56
*** Written on Sat Feb 08, 2025 13:23:47 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

*** SUBCIRCUIT ese3700__nand2 FROM CELL nand2{sch}
.SUBCKT ese3700__nand2 A B Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out A net@1 gnd N L=0.044U W=0.044U
Mnmos@1 net@1 B gnd gnd N L=0.044U W=0.044U
Mpmos@0 vdd B Out vdd P L=0.044U W=0.044U
Mpmos@1 vdd A Out vdd P L=0.044U W=0.044U
.ENDS ese3700__nand2

.global gnd vdd

*** TOP LEVEL CELL: hw2_tranisient{sch}
VVPulse@0 net@30 gnd pulse (0 0.8V 50ps 10ps 10ps 250ps 500ps) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
VV_Generi@1 net@27 gnd DC 0.8 AC 0
VV_Generi@2 net@20 gnd DC 0.8 AC 0
Xnand2@0 MeasureHere1 MeasureHere1 nand2@0_Out ese3700__nand2
Xnand2@1 MeasureHere2 MeasureHere2 nand2@1_Out ese3700__nand2
Xnand2@2 MeasureHere2 MeasureHere2 nand2@2_Out ese3700__nand2
Xnand2@3 MeasureHere1 net@20 MeasureHere2 ese3700__nand2
Xnand2@4 MeasureHere1 net@20 nand2@4_Out ese3700__nand2
Xnand2@5 net@30 net@27 MeasureHere1 ese3700__nand2
.END
