*** SPICE deck for cell hw3_5b{sch} from library ese3700
*** Created on Wed Feb 12, 2025 15:38:37
*** Last revised on Wed Feb 12, 2025 15:58:21
*** Written on Wed Feb 12, 2025 15:58:28 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: hw3_5b{sch}
Mnmos@0 net@0 net@4 gnd gnd N L=0.022U W=0.022U
Mnmos@1 vdd net@0 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@4 net@0 vdd P L=0.022U W=0.022U
VVPulse@0 net@4 gnd pulse (0 0.8V 5ps 0.1ps 1ps 250ps 500ps) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
.END
