*** SPICE deck for cell hw3_6b{sch} from library ese3700
*** Created on Wed Feb 12, 2025 15:01:39
*** Last revised on Wed Feb 12, 2025 15:03:21
*** Written on Wed Feb 12, 2025 15:04:16 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:/Users/garre/ese_3700/22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: hw3_6b{sch}
Mnmos@0 vdd IN OUT gnd N L=0.022U W=0.022U
Mpmos@0 OUT IN gnd vdd P L=0.022U W=0.022U
.END
